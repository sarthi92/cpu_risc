module adder(sum,ain,bin);
output [15:0]sum;
input [15:0]ain,bin;
assign sum=ain+bin;
endmodule
